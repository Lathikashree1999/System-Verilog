interface operation;
  
  logic D;
  logic clk;
  logic rst;
  logic Q;
  
endinterface
