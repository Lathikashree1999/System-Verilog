class transaction;
  
  rand bit D;
  bit clk;
  rand bit rst;
  bit Q;
  
endclass
