interface inter;
  logic a,b,c;
  bit sum,carry;
endinterface
